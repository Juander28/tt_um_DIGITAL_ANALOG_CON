MACRO CON_IV_phvt_nn
  CLASS BLOCK ;
  FOREIGN CON_IV_phvt_nn ;
  ORIGIN -24.640 -6.060 ;
  SIZE 31.440 BY 8.300 ;
  PIN VDD
    ANTENNAGATEAREA 26.000000 ;
    ANTENNADIFFAREA 27.285349 ;
    PORT
      LAYER met1 ;
        RECT 39.515 14.045 40.515 14.165 ;
    END
  END VDD
  PIN GND
    ANTENNAGATEAREA 52.000000 ;
    ANTENNADIFFAREA 16.142099 ;
    PORT
      LAYER met1 ;
        RECT 39.605 6.105 40.605 6.200 ;
    END
  END GND
  PIN N
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER met1 ;
        RECT 41.235 8.750 42.235 8.810 ;
    END
  END N
  PIN P
    ANTENNAGATEAREA 32.000000 ;
    PORT
      LAYER met1 ;
        RECT 41.340 9.350 42.340 9.445 ;
    END
  END P
  PIN VM
    ANTENNAGATEAREA 6.000000 ;
    ANTENNADIFFAREA 1.740000 ;
    PORT
      LAYER met1 ;
        RECT 34.945 9.050 35.945 9.170 ;
    END
  END VM
  OBS
      LAYER nwell ;
        RECT 24.640 9.230 56.080 14.360 ;
      LAYER li1 ;
        RECT 24.685 6.090 56.075 14.175 ;
      LAYER met1 ;
        RECT 24.835 13.765 39.235 14.225 ;
        RECT 40.795 13.765 55.940 14.225 ;
        RECT 24.835 9.725 55.940 13.765 ;
        RECT 24.835 9.450 41.060 9.725 ;
        RECT 24.835 8.770 34.665 9.450 ;
        RECT 36.225 9.090 41.060 9.450 ;
        RECT 36.225 8.770 40.955 9.090 ;
        RECT 42.620 9.070 55.940 9.725 ;
        RECT 24.835 8.470 40.955 8.770 ;
        RECT 42.515 8.470 55.940 9.070 ;
        RECT 24.835 6.480 55.940 8.470 ;
        RECT 24.835 6.060 39.325 6.480 ;
        RECT 40.885 6.060 55.940 6.480 ;
  END
END CON_IV_phvt_nn
END LIBRARY

